class ATM_coverage extends uvm_subscriber;
 
  `uvm_component_utils (ATM_coverage)
  function new(string name = "ATM_coverage");
    super.new(name);
  endfunction
  endclass